// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
// CREATED		"Wed Dec 22 03:05:28 2021"

module tape_64(
	clk,
	rst_n,
	trigger,
	Din,
	keypad,
	pos,
	s,
	tapeData
);


input wire	clk;
input wire	rst_n;
input wire	trigger;
input wire	[1:0] Din;
input wire	[2:0] keypad;
input wire	[5:0] pos;
input wire	[13:0] s;
output wire	[127:0] tapeData;

wire	[127:0] tapeData_ALTERA_SYNTHESIZED;
wire	SYNTHESIZED_WIRE_0;
wire	[1:0] SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_260;
wire	[1:0] SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_5;
wire	[1:0] SYNTHESIZED_WIRE_7;
wire	[1:0] SYNTHESIZED_WIRE_8;
wire	[1:0] SYNTHESIZED_WIRE_9;
wire	[1:0] SYNTHESIZED_WIRE_10;
wire	[1:0] SYNTHESIZED_WIRE_11;
wire	[1:0] SYNTHESIZED_WIRE_12;
wire	[1:0] SYNTHESIZED_WIRE_13;
wire	[1:0] SYNTHESIZED_WIRE_14;
wire	[1:0] SYNTHESIZED_WIRE_15;
wire	[1:0] SYNTHESIZED_WIRE_16;
wire	[1:0] SYNTHESIZED_WIRE_17;
wire	SYNTHESIZED_WIRE_18;
wire	[1:0] SYNTHESIZED_WIRE_20;
wire	[1:0] SYNTHESIZED_WIRE_21;
wire	[1:0] SYNTHESIZED_WIRE_22;
wire	[1:0] SYNTHESIZED_WIRE_23;
wire	[1:0] SYNTHESIZED_WIRE_24;
wire	[1:0] SYNTHESIZED_WIRE_25;
wire	[1:0] SYNTHESIZED_WIRE_26;
wire	[1:0] SYNTHESIZED_WIRE_27;
wire	[1:0] SYNTHESIZED_WIRE_28;
wire	[1:0] SYNTHESIZED_WIRE_29;
wire	[1:0] SYNTHESIZED_WIRE_30;
wire	SYNTHESIZED_WIRE_31;
wire	[1:0] SYNTHESIZED_WIRE_33;
wire	[1:0] SYNTHESIZED_WIRE_34;
wire	[1:0] SYNTHESIZED_WIRE_35;
wire	[1:0] SYNTHESIZED_WIRE_36;
wire	[1:0] SYNTHESIZED_WIRE_37;
wire	[1:0] SYNTHESIZED_WIRE_38;
wire	[1:0] SYNTHESIZED_WIRE_39;
wire	[1:0] SYNTHESIZED_WIRE_40;
wire	[1:0] SYNTHESIZED_WIRE_41;
wire	[1:0] SYNTHESIZED_WIRE_42;
wire	[1:0] SYNTHESIZED_WIRE_43;
wire	SYNTHESIZED_WIRE_44;
wire	[1:0] SYNTHESIZED_WIRE_46;
wire	[1:0] SYNTHESIZED_WIRE_47;
wire	SYNTHESIZED_WIRE_48;
wire	SYNTHESIZED_WIRE_49;
wire	[1:0] SYNTHESIZED_WIRE_51;
wire	SYNTHESIZED_WIRE_52;
wire	[1:0] SYNTHESIZED_WIRE_54;
wire	SYNTHESIZED_WIRE_55;
wire	[1:0] SYNTHESIZED_WIRE_57;
wire	SYNTHESIZED_WIRE_58;
wire	[1:0] SYNTHESIZED_WIRE_60;
wire	SYNTHESIZED_WIRE_61;
wire	[1:0] SYNTHESIZED_WIRE_63;
wire	SYNTHESIZED_WIRE_64;
wire	[1:0] SYNTHESIZED_WIRE_66;
wire	SYNTHESIZED_WIRE_67;
wire	[1:0] SYNTHESIZED_WIRE_69;
wire	SYNTHESIZED_WIRE_70;
wire	[1:0] SYNTHESIZED_WIRE_72;
wire	SYNTHESIZED_WIRE_73;
wire	[1:0] SYNTHESIZED_WIRE_75;
wire	SYNTHESIZED_WIRE_76;
wire	[1:0] SYNTHESIZED_WIRE_78;
wire	SYNTHESIZED_WIRE_79;
wire	[1:0] SYNTHESIZED_WIRE_81;
wire	SYNTHESIZED_WIRE_82;
wire	[1:0] SYNTHESIZED_WIRE_84;
wire	SYNTHESIZED_WIRE_85;
wire	[1:0] SYNTHESIZED_WIRE_87;
wire	SYNTHESIZED_WIRE_88;
wire	[1:0] SYNTHESIZED_WIRE_90;
wire	SYNTHESIZED_WIRE_91;
wire	[1:0] SYNTHESIZED_WIRE_93;
wire	SYNTHESIZED_WIRE_94;
wire	[1:0] SYNTHESIZED_WIRE_96;
wire	SYNTHESIZED_WIRE_97;
wire	[1:0] SYNTHESIZED_WIRE_99;
wire	SYNTHESIZED_WIRE_100;
wire	[1:0] SYNTHESIZED_WIRE_102;
wire	SYNTHESIZED_WIRE_103;
wire	[1:0] SYNTHESIZED_WIRE_105;
wire	SYNTHESIZED_WIRE_106;
wire	[1:0] SYNTHESIZED_WIRE_108;
wire	SYNTHESIZED_WIRE_109;
wire	[1:0] SYNTHESIZED_WIRE_111;
wire	SYNTHESIZED_WIRE_112;
wire	[1:0] SYNTHESIZED_WIRE_114;
wire	SYNTHESIZED_WIRE_115;
wire	[1:0] SYNTHESIZED_WIRE_117;
wire	SYNTHESIZED_WIRE_118;
wire	[1:0] SYNTHESIZED_WIRE_120;
wire	SYNTHESIZED_WIRE_121;
wire	[1:0] SYNTHESIZED_WIRE_123;
wire	SYNTHESIZED_WIRE_124;
wire	[1:0] SYNTHESIZED_WIRE_126;
wire	SYNTHESIZED_WIRE_127;
wire	[1:0] SYNTHESIZED_WIRE_129;
wire	SYNTHESIZED_WIRE_130;
wire	[1:0] SYNTHESIZED_WIRE_132;
wire	SYNTHESIZED_WIRE_133;
wire	[1:0] SYNTHESIZED_WIRE_135;
wire	SYNTHESIZED_WIRE_136;
wire	[1:0] SYNTHESIZED_WIRE_138;
wire	SYNTHESIZED_WIRE_139;
wire	[1:0] SYNTHESIZED_WIRE_141;
wire	SYNTHESIZED_WIRE_142;
wire	[1:0] SYNTHESIZED_WIRE_144;
wire	SYNTHESIZED_WIRE_145;
wire	[1:0] SYNTHESIZED_WIRE_147;
wire	SYNTHESIZED_WIRE_148;
wire	[1:0] SYNTHESIZED_WIRE_150;
wire	SYNTHESIZED_WIRE_151;
wire	[1:0] SYNTHESIZED_WIRE_153;
wire	SYNTHESIZED_WIRE_154;
wire	[1:0] SYNTHESIZED_WIRE_156;
wire	SYNTHESIZED_WIRE_157;
wire	[1:0] SYNTHESIZED_WIRE_159;
wire	SYNTHESIZED_WIRE_160;
wire	[1:0] SYNTHESIZED_WIRE_162;
wire	SYNTHESIZED_WIRE_163;
wire	[1:0] SYNTHESIZED_WIRE_165;
wire	SYNTHESIZED_WIRE_166;
wire	[1:0] SYNTHESIZED_WIRE_168;
wire	SYNTHESIZED_WIRE_169;
wire	[1:0] SYNTHESIZED_WIRE_171;
wire	SYNTHESIZED_WIRE_172;
wire	[1:0] SYNTHESIZED_WIRE_174;
wire	SYNTHESIZED_WIRE_175;
wire	[1:0] SYNTHESIZED_WIRE_177;
wire	SYNTHESIZED_WIRE_178;
wire	[1:0] SYNTHESIZED_WIRE_180;
wire	SYNTHESIZED_WIRE_181;
wire	[1:0] SYNTHESIZED_WIRE_183;
wire	SYNTHESIZED_WIRE_184;
wire	[1:0] SYNTHESIZED_WIRE_186;
wire	SYNTHESIZED_WIRE_187;
wire	[1:0] SYNTHESIZED_WIRE_189;
wire	SYNTHESIZED_WIRE_190;
wire	[1:0] SYNTHESIZED_WIRE_192;
wire	SYNTHESIZED_WIRE_193;
wire	[1:0] SYNTHESIZED_WIRE_195;
wire	SYNTHESIZED_WIRE_196;
wire	[1:0] SYNTHESIZED_WIRE_198;
wire	SYNTHESIZED_WIRE_199;
wire	[1:0] SYNTHESIZED_WIRE_201;
wire	SYNTHESIZED_WIRE_202;
wire	[1:0] SYNTHESIZED_WIRE_204;
wire	SYNTHESIZED_WIRE_205;
wire	[1:0] SYNTHESIZED_WIRE_207;
wire	SYNTHESIZED_WIRE_208;
wire	[1:0] SYNTHESIZED_WIRE_210;
wire	SYNTHESIZED_WIRE_211;
wire	[1:0] SYNTHESIZED_WIRE_213;
wire	SYNTHESIZED_WIRE_214;
wire	[1:0] SYNTHESIZED_WIRE_216;
wire	SYNTHESIZED_WIRE_217;
wire	[1:0] SYNTHESIZED_WIRE_218;
wire	[1:0] SYNTHESIZED_WIRE_219;
wire	[1:0] SYNTHESIZED_WIRE_220;
wire	SYNTHESIZED_WIRE_221;
wire	[1:0] SYNTHESIZED_WIRE_223;
wire	[1:0] SYNTHESIZED_WIRE_224;
wire	[1:0] SYNTHESIZED_WIRE_225;
wire	[1:0] SYNTHESIZED_WIRE_226;
wire	[1:0] SYNTHESIZED_WIRE_227;
wire	[1:0] SYNTHESIZED_WIRE_228;
wire	[1:0] SYNTHESIZED_WIRE_229;
wire	[1:0] SYNTHESIZED_WIRE_230;
wire	[1:0] SYNTHESIZED_WIRE_231;
wire	[1:0] SYNTHESIZED_WIRE_232;
wire	[1:0] SYNTHESIZED_WIRE_233;
wire	SYNTHESIZED_WIRE_234;
wire	[1:0] SYNTHESIZED_WIRE_236;
wire	[1:0] SYNTHESIZED_WIRE_237;
wire	[1:0] SYNTHESIZED_WIRE_238;
wire	[1:0] SYNTHESIZED_WIRE_239;
wire	[1:0] SYNTHESIZED_WIRE_240;
wire	[1:0] SYNTHESIZED_WIRE_241;
wire	[1:0] SYNTHESIZED_WIRE_242;
wire	[1:0] SYNTHESIZED_WIRE_243;
wire	[1:0] SYNTHESIZED_WIRE_244;
wire	[1:0] SYNTHESIZED_WIRE_245;
wire	[1:0] SYNTHESIZED_WIRE_246;
wire	SYNTHESIZED_WIRE_247;
wire	[1:0] SYNTHESIZED_WIRE_249;
wire	[1:0] SYNTHESIZED_WIRE_250;
wire	[1:0] SYNTHESIZED_WIRE_251;
wire	[1:0] SYNTHESIZED_WIRE_252;
wire	[1:0] SYNTHESIZED_WIRE_253;
wire	[1:0] SYNTHESIZED_WIRE_254;
wire	[1:0] SYNTHESIZED_WIRE_255;
wire	[1:0] SYNTHESIZED_WIRE_256;
wire	[1:0] SYNTHESIZED_WIRE_257;
wire	[1:0] SYNTHESIZED_WIRE_258;
wire	[1:0] SYNTHESIZED_WIRE_259;




assign	SYNTHESIZED_WIRE_260 = SYNTHESIZED_WIRE_0 & rst_n;


Mux2bit2x1	b2v_dinmux(
	.sel(s[1]),
	.Din0(Din),
	.Din1(keypad[1:0]),
	.Dout(SYNTHESIZED_WIRE_1));


demux_1x64_2bit	b2v_inst(
	.Din(SYNTHESIZED_WIRE_1),
	.sel(pos),
	.Dout_0_(SYNTHESIZED_WIRE_4),
	.Dout_10_(SYNTHESIZED_WIRE_20),
	.Dout_11_(SYNTHESIZED_WIRE_33),
	.Dout_12_(SYNTHESIZED_WIRE_46),
	.Dout_13_(SYNTHESIZED_WIRE_51),
	.Dout_14_(SYNTHESIZED_WIRE_54),
	.Dout_15_(SYNTHESIZED_WIRE_57),
	.Dout_16_(SYNTHESIZED_WIRE_60),
	.Dout_17_(SYNTHESIZED_WIRE_63),
	.Dout_18_(SYNTHESIZED_WIRE_66),
	.Dout_19_(SYNTHESIZED_WIRE_72),
	.Dout_1_(SYNTHESIZED_WIRE_69),
	.Dout_20_(SYNTHESIZED_WIRE_75),
	.Dout_21_(SYNTHESIZED_WIRE_78),
	.Dout_22_(SYNTHESIZED_WIRE_81),
	.Dout_23_(SYNTHESIZED_WIRE_84),
	.Dout_24_(SYNTHESIZED_WIRE_87),
	.Dout_25_(SYNTHESIZED_WIRE_90),
	.Dout_26_(SYNTHESIZED_WIRE_93),
	.Dout_27_(SYNTHESIZED_WIRE_96),
	.Dout_28_(SYNTHESIZED_WIRE_99),
	.Dout_29_(SYNTHESIZED_WIRE_105),
	.Dout_2_(SYNTHESIZED_WIRE_102),
	.Dout_30_(SYNTHESIZED_WIRE_108),
	.Dout_31_(SYNTHESIZED_WIRE_111),
	.Dout_32_(SYNTHESIZED_WIRE_114),
	.Dout_33_(SYNTHESIZED_WIRE_117),
	.Dout_34_(SYNTHESIZED_WIRE_120),
	.Dout_35_(SYNTHESIZED_WIRE_123),
	.Dout_36_(SYNTHESIZED_WIRE_126),
	.Dout_37_(SYNTHESIZED_WIRE_129),
	.Dout_38_(SYNTHESIZED_WIRE_132),
	.Dout_39_(SYNTHESIZED_WIRE_138),
	.Dout_3_(SYNTHESIZED_WIRE_135),
	.Dout_40_(SYNTHESIZED_WIRE_141),
	.Dout_41_(SYNTHESIZED_WIRE_144),
	.Dout_42_(SYNTHESIZED_WIRE_147),
	.Dout_43_(SYNTHESIZED_WIRE_150),
	.Dout_44_(SYNTHESIZED_WIRE_153),
	.Dout_45_(SYNTHESIZED_WIRE_156),
	.Dout_46_(SYNTHESIZED_WIRE_159),
	.Dout_47_(SYNTHESIZED_WIRE_162),
	.Dout_48_(SYNTHESIZED_WIRE_165),
	.Dout_49_(SYNTHESIZED_WIRE_171),
	.Dout_4_(SYNTHESIZED_WIRE_168),
	.Dout_50_(SYNTHESIZED_WIRE_174),
	.Dout_51_(SYNTHESIZED_WIRE_177),
	.Dout_52_(SYNTHESIZED_WIRE_180),
	.Dout_53_(SYNTHESIZED_WIRE_183),
	.Dout_54_(SYNTHESIZED_WIRE_186),
	.Dout_55_(SYNTHESIZED_WIRE_189),
	.Dout_56_(SYNTHESIZED_WIRE_192),
	.Dout_57_(SYNTHESIZED_WIRE_195),
	.Dout_58_(SYNTHESIZED_WIRE_198),
	.Dout_59_(SYNTHESIZED_WIRE_204),
	.Dout_5_(SYNTHESIZED_WIRE_201),
	.Dout_60_(SYNTHESIZED_WIRE_207),
	.Dout_61_(SYNTHESIZED_WIRE_210),
	.Dout_62_(SYNTHESIZED_WIRE_213),
	.Dout_63_(SYNTHESIZED_WIRE_216),
	.Dout_6_(SYNTHESIZED_WIRE_223),
	.Dout_7_(SYNTHESIZED_WIRE_236),
	.Dout_8_(SYNTHESIZED_WIRE_249),
	.Dout_9_(SYNTHESIZED_WIRE_7));


reg_2bit	b2v_inst1(
	.Ce(SYNTHESIZED_WIRE_2),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_4),
	.Dout(SYNTHESIZED_WIRE_218));


reg_2bit	b2v_inst10(
	.Ce(SYNTHESIZED_WIRE_5),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_7),
	.Dout(SYNTHESIZED_WIRE_230));


cvt_2x1_1x2	b2v_inst100(
	.Din(SYNTHESIZED_WIRE_8),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[66]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[67]));


cvt_2x1_1x2	b2v_inst101(
	.Din(SYNTHESIZED_WIRE_9),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[68]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[69]));


cvt_2x1_1x2	b2v_inst102(
	.Din(SYNTHESIZED_WIRE_10),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[70]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[71]));


cvt_2x1_1x2	b2v_inst103(
	.Din(SYNTHESIZED_WIRE_11),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[72]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[73]));


cvt_2x1_1x2	b2v_inst104(
	.Din(SYNTHESIZED_WIRE_12),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[74]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[75]));


cvt_2x1_1x2	b2v_inst105(
	.Din(SYNTHESIZED_WIRE_13),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[76]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[77]));


cvt_2x1_1x2	b2v_inst106(
	.Din(SYNTHESIZED_WIRE_14),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[78]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[79]));


cvt_2x1_1x2	b2v_inst107(
	.Din(SYNTHESIZED_WIRE_15),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[80]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[81]));


cvt_2x1_1x2	b2v_inst108(
	.Din(SYNTHESIZED_WIRE_16),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[82]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[83]));


cvt_2x1_1x2	b2v_inst109(
	.Din(SYNTHESIZED_WIRE_17),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[84]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[85]));


reg_2bit	b2v_inst11(
	.Ce(SYNTHESIZED_WIRE_18),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_20),
	.Dout(SYNTHESIZED_WIRE_231));


cvt_2x1_1x2	b2v_inst110(
	.Din(SYNTHESIZED_WIRE_21),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[86]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[87]));


cvt_2x1_1x2	b2v_inst111(
	.Din(SYNTHESIZED_WIRE_22),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[88]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[89]));


cvt_2x1_1x2	b2v_inst112(
	.Din(SYNTHESIZED_WIRE_23),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[90]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[91]));


cvt_2x1_1x2	b2v_inst113(
	.Din(SYNTHESIZED_WIRE_24),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[92]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[93]));


cvt_2x1_1x2	b2v_inst114(
	.Din(SYNTHESIZED_WIRE_25),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[94]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[95]));


cvt_2x1_1x2	b2v_inst115(
	.Din(SYNTHESIZED_WIRE_26),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[96]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[97]));


cvt_2x1_1x2	b2v_inst116(
	.Din(SYNTHESIZED_WIRE_27),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[98]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[99]));


cvt_2x1_1x2	b2v_inst117(
	.Din(SYNTHESIZED_WIRE_28),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[100]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[101]));


cvt_2x1_1x2	b2v_inst118(
	.Din(SYNTHESIZED_WIRE_29),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[102]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[103]));


cvt_2x1_1x2	b2v_inst119(
	.Din(SYNTHESIZED_WIRE_30),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[104]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[105]));


reg_2bit	b2v_inst12(
	.Ce(SYNTHESIZED_WIRE_31),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_33),
	.Dout(SYNTHESIZED_WIRE_232));


cvt_2x1_1x2	b2v_inst120(
	.Din(SYNTHESIZED_WIRE_34),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[106]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[107]));


cvt_2x1_1x2	b2v_inst121(
	.Din(SYNTHESIZED_WIRE_35),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[108]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[109]));


cvt_2x1_1x2	b2v_inst122(
	.Din(SYNTHESIZED_WIRE_36),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[110]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[111]));


cvt_2x1_1x2	b2v_inst123(
	.Din(SYNTHESIZED_WIRE_37),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[112]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[113]));


cvt_2x1_1x2	b2v_inst124(
	.Din(SYNTHESIZED_WIRE_38),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[114]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[115]));


cvt_2x1_1x2	b2v_inst125(
	.Din(SYNTHESIZED_WIRE_39),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[116]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[117]));


cvt_2x1_1x2	b2v_inst126(
	.Din(SYNTHESIZED_WIRE_40),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[118]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[119]));


cvt_2x1_1x2	b2v_inst127(
	.Din(SYNTHESIZED_WIRE_41),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[120]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[121]));


cvt_2x1_1x2	b2v_inst128(
	.Din(SYNTHESIZED_WIRE_42),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[122]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[123]));


cvt_2x1_1x2	b2v_inst129(
	.Din(SYNTHESIZED_WIRE_43),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[124]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[125]));


reg_2bit	b2v_inst13(
	.Ce(SYNTHESIZED_WIRE_44),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_46),
	.Dout(SYNTHESIZED_WIRE_233));


cvt_2x1_1x2	b2v_inst130(
	.Din(SYNTHESIZED_WIRE_47),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[126]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[127]));

assign	SYNTHESIZED_WIRE_217 = s[10] | SYNTHESIZED_WIRE_48;


reg_2bit	b2v_inst14(
	.Ce(SYNTHESIZED_WIRE_49),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_51),
	.Dout(SYNTHESIZED_WIRE_237));


reg_2bit	b2v_inst15(
	.Ce(SYNTHESIZED_WIRE_52),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_54),
	.Dout(SYNTHESIZED_WIRE_238));


reg_2bit	b2v_inst16(
	.Ce(SYNTHESIZED_WIRE_55),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_57),
	.Dout(SYNTHESIZED_WIRE_239));


reg_2bit	b2v_inst17(
	.Ce(SYNTHESIZED_WIRE_58),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_60),
	.Dout(SYNTHESIZED_WIRE_240));


reg_2bit	b2v_inst18(
	.Ce(SYNTHESIZED_WIRE_61),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_63),
	.Dout(SYNTHESIZED_WIRE_241));


reg_2bit	b2v_inst19(
	.Ce(SYNTHESIZED_WIRE_64),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_66),
	.Dout(SYNTHESIZED_WIRE_242));


reg_2bit	b2v_inst2(
	.Ce(SYNTHESIZED_WIRE_67),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_69),
	.Dout(SYNTHESIZED_WIRE_219));


reg_2bit	b2v_inst20(
	.Ce(SYNTHESIZED_WIRE_70),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_72),
	.Dout(SYNTHESIZED_WIRE_243));


reg_2bit	b2v_inst21(
	.Ce(SYNTHESIZED_WIRE_73),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_75),
	.Dout(SYNTHESIZED_WIRE_244));


reg_2bit	b2v_inst22(
	.Ce(SYNTHESIZED_WIRE_76),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_78),
	.Dout(SYNTHESIZED_WIRE_245));


reg_2bit	b2v_inst23(
	.Ce(SYNTHESIZED_WIRE_79),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_81),
	.Dout(SYNTHESIZED_WIRE_246));


reg_2bit	b2v_inst24(
	.Ce(SYNTHESIZED_WIRE_82),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_84),
	.Dout(SYNTHESIZED_WIRE_250));


reg_2bit	b2v_inst25(
	.Ce(SYNTHESIZED_WIRE_85),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_87),
	.Dout(SYNTHESIZED_WIRE_251));


reg_2bit	b2v_inst26(
	.Ce(SYNTHESIZED_WIRE_88),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_90),
	.Dout(SYNTHESIZED_WIRE_252));


reg_2bit	b2v_inst27(
	.Ce(SYNTHESIZED_WIRE_91),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_93),
	.Dout(SYNTHESIZED_WIRE_253));


reg_2bit	b2v_inst28(
	.Ce(SYNTHESIZED_WIRE_94),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_96),
	.Dout(SYNTHESIZED_WIRE_254));


reg_2bit	b2v_inst29(
	.Ce(SYNTHESIZED_WIRE_97),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_99),
	.Dout(SYNTHESIZED_WIRE_255));


reg_2bit	b2v_inst3(
	.Ce(SYNTHESIZED_WIRE_100),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_102),
	.Dout(SYNTHESIZED_WIRE_220));


reg_2bit	b2v_inst30(
	.Ce(SYNTHESIZED_WIRE_103),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_105),
	.Dout(SYNTHESIZED_WIRE_256));


reg_2bit	b2v_inst31(
	.Ce(SYNTHESIZED_WIRE_106),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_108),
	.Dout(SYNTHESIZED_WIRE_257));


reg_2bit	b2v_inst32(
	.Ce(SYNTHESIZED_WIRE_109),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_111),
	.Dout(SYNTHESIZED_WIRE_258));


reg_2bit	b2v_inst33(
	.Ce(SYNTHESIZED_WIRE_112),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_114),
	.Dout(SYNTHESIZED_WIRE_259));


reg_2bit	b2v_inst34(
	.Ce(SYNTHESIZED_WIRE_115),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_117),
	.Dout(SYNTHESIZED_WIRE_8));


reg_2bit	b2v_inst35(
	.Ce(SYNTHESIZED_WIRE_118),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_120),
	.Dout(SYNTHESIZED_WIRE_9));


reg_2bit	b2v_inst36(
	.Ce(SYNTHESIZED_WIRE_121),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_123),
	.Dout(SYNTHESIZED_WIRE_10));


reg_2bit	b2v_inst37(
	.Ce(SYNTHESIZED_WIRE_124),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_126),
	.Dout(SYNTHESIZED_WIRE_11));


reg_2bit	b2v_inst38(
	.Ce(SYNTHESIZED_WIRE_127),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_129),
	.Dout(SYNTHESIZED_WIRE_12));


reg_2bit	b2v_inst39(
	.Ce(SYNTHESIZED_WIRE_130),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_132),
	.Dout(SYNTHESIZED_WIRE_13));


reg_2bit	b2v_inst4(
	.Ce(SYNTHESIZED_WIRE_133),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_135),
	.Dout(SYNTHESIZED_WIRE_224));


reg_2bit	b2v_inst40(
	.Ce(SYNTHESIZED_WIRE_136),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_138),
	.Dout(SYNTHESIZED_WIRE_14));


reg_2bit	b2v_inst41(
	.Ce(SYNTHESIZED_WIRE_139),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_141),
	.Dout(SYNTHESIZED_WIRE_15));


reg_2bit	b2v_inst42(
	.Ce(SYNTHESIZED_WIRE_142),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_144),
	.Dout(SYNTHESIZED_WIRE_16));


reg_2bit	b2v_inst43(
	.Ce(SYNTHESIZED_WIRE_145),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_147),
	.Dout(SYNTHESIZED_WIRE_17));


reg_2bit	b2v_inst44(
	.Ce(SYNTHESIZED_WIRE_148),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_150),
	.Dout(SYNTHESIZED_WIRE_21));


reg_2bit	b2v_inst45(
	.Ce(SYNTHESIZED_WIRE_151),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_153),
	.Dout(SYNTHESIZED_WIRE_22));


reg_2bit	b2v_inst46(
	.Ce(SYNTHESIZED_WIRE_154),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_156),
	.Dout(SYNTHESIZED_WIRE_23));


reg_2bit	b2v_inst47(
	.Ce(SYNTHESIZED_WIRE_157),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_159),
	.Dout(SYNTHESIZED_WIRE_24));


reg_2bit	b2v_inst48(
	.Ce(SYNTHESIZED_WIRE_160),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_162),
	.Dout(SYNTHESIZED_WIRE_25));


reg_2bit	b2v_inst49(
	.Ce(SYNTHESIZED_WIRE_163),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_165),
	.Dout(SYNTHESIZED_WIRE_26));


reg_2bit	b2v_inst5(
	.Ce(SYNTHESIZED_WIRE_166),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_168),
	.Dout(SYNTHESIZED_WIRE_225));


reg_2bit	b2v_inst50(
	.Ce(SYNTHESIZED_WIRE_169),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_171),
	.Dout(SYNTHESIZED_WIRE_27));


reg_2bit	b2v_inst51(
	.Ce(SYNTHESIZED_WIRE_172),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_174),
	.Dout(SYNTHESIZED_WIRE_28));


reg_2bit	b2v_inst52(
	.Ce(SYNTHESIZED_WIRE_175),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_177),
	.Dout(SYNTHESIZED_WIRE_29));


reg_2bit	b2v_inst53(
	.Ce(SYNTHESIZED_WIRE_178),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_180),
	.Dout(SYNTHESIZED_WIRE_30));


reg_2bit	b2v_inst54(
	.Ce(SYNTHESIZED_WIRE_181),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_183),
	.Dout(SYNTHESIZED_WIRE_34));


reg_2bit	b2v_inst55(
	.Ce(SYNTHESIZED_WIRE_184),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_186),
	.Dout(SYNTHESIZED_WIRE_35));


reg_2bit	b2v_inst56(
	.Ce(SYNTHESIZED_WIRE_187),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_189),
	.Dout(SYNTHESIZED_WIRE_36));


reg_2bit	b2v_inst57(
	.Ce(SYNTHESIZED_WIRE_190),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_192),
	.Dout(SYNTHESIZED_WIRE_37));


reg_2bit	b2v_inst58(
	.Ce(SYNTHESIZED_WIRE_193),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_195),
	.Dout(SYNTHESIZED_WIRE_38));


reg_2bit	b2v_inst59(
	.Ce(SYNTHESIZED_WIRE_196),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_198),
	.Dout(SYNTHESIZED_WIRE_39));


reg_2bit	b2v_inst6(
	.Ce(SYNTHESIZED_WIRE_199),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_201),
	.Dout(SYNTHESIZED_WIRE_226));


reg_2bit	b2v_inst60(
	.Ce(SYNTHESIZED_WIRE_202),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_204),
	.Dout(SYNTHESIZED_WIRE_40));


reg_2bit	b2v_inst61(
	.Ce(SYNTHESIZED_WIRE_205),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_207),
	.Dout(SYNTHESIZED_WIRE_41));


reg_2bit	b2v_inst62(
	.Ce(SYNTHESIZED_WIRE_208),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_210),
	.Dout(SYNTHESIZED_WIRE_42));


reg_2bit	b2v_inst63(
	.Ce(SYNTHESIZED_WIRE_211),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_213),
	.Dout(SYNTHESIZED_WIRE_43));


reg_2bit	b2v_inst64(
	.Ce(SYNTHESIZED_WIRE_214),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_216),
	.Dout(SYNTHESIZED_WIRE_47));


demux_1x64	b2v_inst65(
	.Din(SYNTHESIZED_WIRE_217),
	.sel(pos),
	.Dout_63(SYNTHESIZED_WIRE_214),
	.Dout_62(SYNTHESIZED_WIRE_211),
	.Dout_61(SYNTHESIZED_WIRE_208),
	.Dout_60(SYNTHESIZED_WIRE_205),
	.Dout_59(SYNTHESIZED_WIRE_202),
	.Dout_58(SYNTHESIZED_WIRE_196),
	.Dout_57(SYNTHESIZED_WIRE_193),
	.Dout_56(SYNTHESIZED_WIRE_190),
	.Dout_55(SYNTHESIZED_WIRE_187),
	.Dout_54(SYNTHESIZED_WIRE_184),
	.Dout_53(SYNTHESIZED_WIRE_181),
	.Dout_52(SYNTHESIZED_WIRE_178),
	.Dout_51(SYNTHESIZED_WIRE_175),
	.Dout_50(SYNTHESIZED_WIRE_172),
	.Dout_49(SYNTHESIZED_WIRE_169),
	.Dout_48(SYNTHESIZED_WIRE_163),
	.Dout_47(SYNTHESIZED_WIRE_160),
	.Dout_46(SYNTHESIZED_WIRE_157),
	.Dout_45(SYNTHESIZED_WIRE_154),
	.Dout_44(SYNTHESIZED_WIRE_151),
	.Dout_43(SYNTHESIZED_WIRE_148),
	.Dout_42(SYNTHESIZED_WIRE_145),
	.Dout_41(SYNTHESIZED_WIRE_142),
	.Dout_40(SYNTHESIZED_WIRE_139),
	.Dout_39(SYNTHESIZED_WIRE_136),
	.Dout_38(SYNTHESIZED_WIRE_130),
	.Dout_37(SYNTHESIZED_WIRE_127),
	.Dout_36(SYNTHESIZED_WIRE_124),
	.Dout_35(SYNTHESIZED_WIRE_121),
	.Dout_34(SYNTHESIZED_WIRE_118),
	.Dout_33(SYNTHESIZED_WIRE_115),
	.Dout_32(SYNTHESIZED_WIRE_112),
	.Dout_31(SYNTHESIZED_WIRE_109),
	.Dout_30(SYNTHESIZED_WIRE_106),
	.Dout_29(SYNTHESIZED_WIRE_103),
	.Dout_28(SYNTHESIZED_WIRE_97),
	.Dout_27(SYNTHESIZED_WIRE_94),
	.Dout_26(SYNTHESIZED_WIRE_91),
	.Dout_25(SYNTHESIZED_WIRE_88),
	.Dout_24(SYNTHESIZED_WIRE_85),
	.Dout_23(SYNTHESIZED_WIRE_82),
	.Dout_22(SYNTHESIZED_WIRE_79),
	.Dout_21(SYNTHESIZED_WIRE_76),
	.Dout_20(SYNTHESIZED_WIRE_73),
	.Dout_19(SYNTHESIZED_WIRE_70),
	.Dout_18(SYNTHESIZED_WIRE_64),
	.Dout_17(SYNTHESIZED_WIRE_61),
	.Dout_16(SYNTHESIZED_WIRE_58),
	.Dout_15(SYNTHESIZED_WIRE_55),
	.Dout_14(SYNTHESIZED_WIRE_52),
	.Dout_13(SYNTHESIZED_WIRE_49),
	.Dout_12(SYNTHESIZED_WIRE_44),
	.Dout_11(SYNTHESIZED_WIRE_31),
	.Dout_10(SYNTHESIZED_WIRE_18),
	.Dout_9(SYNTHESIZED_WIRE_5),
	.Dout_8(SYNTHESIZED_WIRE_247),
	.Dout_7(SYNTHESIZED_WIRE_234),
	.Dout_6(SYNTHESIZED_WIRE_221),
	.Dout_5(SYNTHESIZED_WIRE_199),
	.Dout_4(SYNTHESIZED_WIRE_166),
	.Dout_3(SYNTHESIZED_WIRE_133),
	.Dout_2(SYNTHESIZED_WIRE_100),
	.Dout_1(SYNTHESIZED_WIRE_67),
	.Dout_0(SYNTHESIZED_WIRE_2));

assign	SYNTHESIZED_WIRE_48 = trigger & s[1];


cvt_2x1_1x2	b2v_inst67(
	.Din(SYNTHESIZED_WIRE_218),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[0]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[1]));


cvt_2x1_1x2	b2v_inst68(
	.Din(SYNTHESIZED_WIRE_219),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[2]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[3]));


cvt_2x1_1x2	b2v_inst69(
	.Din(SYNTHESIZED_WIRE_220),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[4]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[5]));


reg_2bit	b2v_inst7(
	.Ce(SYNTHESIZED_WIRE_221),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_223),
	.Dout(SYNTHESIZED_WIRE_227));


cvt_2x1_1x2	b2v_inst70(
	.Din(SYNTHESIZED_WIRE_224),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[6]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[7]));


cvt_2x1_1x2	b2v_inst71(
	.Din(SYNTHESIZED_WIRE_225),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[8]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[9]));


cvt_2x1_1x2	b2v_inst72(
	.Din(SYNTHESIZED_WIRE_226),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[10]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[11]));


cvt_2x1_1x2	b2v_inst73(
	.Din(SYNTHESIZED_WIRE_227),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[12]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[13]));


cvt_2x1_1x2	b2v_inst74(
	.Din(SYNTHESIZED_WIRE_228),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[14]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[15]));


cvt_2x1_1x2	b2v_inst75(
	.Din(SYNTHESIZED_WIRE_229),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[16]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[17]));


cvt_2x1_1x2	b2v_inst76(
	.Din(SYNTHESIZED_WIRE_230),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[18]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[19]));


cvt_2x1_1x2	b2v_inst77(
	.Din(SYNTHESIZED_WIRE_231),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[20]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[21]));


cvt_2x1_1x2	b2v_inst78(
	.Din(SYNTHESIZED_WIRE_232),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[22]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[23]));


cvt_2x1_1x2	b2v_inst79(
	.Din(SYNTHESIZED_WIRE_233),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[24]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[25]));


reg_2bit	b2v_inst8(
	.Ce(SYNTHESIZED_WIRE_234),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_236),
	.Dout(SYNTHESIZED_WIRE_228));


cvt_2x1_1x2	b2v_inst80(
	.Din(SYNTHESIZED_WIRE_237),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[26]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[27]));


cvt_2x1_1x2	b2v_inst81(
	.Din(SYNTHESIZED_WIRE_238),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[28]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[29]));


cvt_2x1_1x2	b2v_inst82(
	.Din(SYNTHESIZED_WIRE_239),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[30]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[31]));


cvt_2x1_1x2	b2v_inst83(
	.Din(SYNTHESIZED_WIRE_240),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[32]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[33]));


cvt_2x1_1x2	b2v_inst84(
	.Din(SYNTHESIZED_WIRE_241),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[34]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[35]));


cvt_2x1_1x2	b2v_inst85(
	.Din(SYNTHESIZED_WIRE_242),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[36]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[37]));


cvt_2x1_1x2	b2v_inst86(
	.Din(SYNTHESIZED_WIRE_243),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[38]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[39]));


cvt_2x1_1x2	b2v_inst87(
	.Din(SYNTHESIZED_WIRE_244),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[40]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[41]));


cvt_2x1_1x2	b2v_inst88(
	.Din(SYNTHESIZED_WIRE_245),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[42]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[43]));


cvt_2x1_1x2	b2v_inst89(
	.Din(SYNTHESIZED_WIRE_246),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[44]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[45]));


reg_2bit	b2v_inst9(
	.Ce(SYNTHESIZED_WIRE_247),
	.clk(clk),
	.rst_n(SYNTHESIZED_WIRE_260),
	.Din(SYNTHESIZED_WIRE_249),
	.Dout(SYNTHESIZED_WIRE_229));


cvt_2x1_1x2	b2v_inst90(
	.Din(SYNTHESIZED_WIRE_250),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[46]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[47]));


cvt_2x1_1x2	b2v_inst91(
	.Din(SYNTHESIZED_WIRE_251),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[48]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[49]));


cvt_2x1_1x2	b2v_inst92(
	.Din(SYNTHESIZED_WIRE_252),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[50]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[51]));


cvt_2x1_1x2	b2v_inst93(
	.Din(SYNTHESIZED_WIRE_253),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[52]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[53]));


cvt_2x1_1x2	b2v_inst94(
	.Din(SYNTHESIZED_WIRE_254),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[54]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[55]));


cvt_2x1_1x2	b2v_inst95(
	.Din(SYNTHESIZED_WIRE_255),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[56]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[57]));


cvt_2x1_1x2	b2v_inst96(
	.Din(SYNTHESIZED_WIRE_256),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[58]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[59]));


cvt_2x1_1x2	b2v_inst97(
	.Din(SYNTHESIZED_WIRE_257),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[60]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[61]));


cvt_2x1_1x2	b2v_inst98(
	.Din(SYNTHESIZED_WIRE_258),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[62]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[63]));


cvt_2x1_1x2	b2v_inst99(
	.Din(SYNTHESIZED_WIRE_259),
	.Dout0(tapeData_ALTERA_SYNTHESIZED[64]),
	.Dout1(tapeData_ALTERA_SYNTHESIZED[65]));

assign	SYNTHESIZED_WIRE_0 =  ~s[13];

assign	tapeData = tapeData_ALTERA_SYNTHESIZED;

endmodule
