// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
// CREATED		"Tue Dec 21 11:58:26 2021"

module tapeSymbolFinder(
	sel,
	tapeData,
	tapeSymbol
);


input wire	[5:0] sel;
input wire	[127:0] tapeData;
output wire	[1:0] tapeSymbol;

wire	[1:0] SYNTHESIZED_WIRE_0;
wire	[1:0] SYNTHESIZED_WIRE_1;
wire	[1:0] SYNTHESIZED_WIRE_2;
wire	[1:0] SYNTHESIZED_WIRE_3;
wire	[1:0] SYNTHESIZED_WIRE_4;
wire	[1:0] SYNTHESIZED_WIRE_5;
wire	[1:0] SYNTHESIZED_WIRE_6;
wire	[1:0] SYNTHESIZED_WIRE_7;
wire	[1:0] SYNTHESIZED_WIRE_8;
wire	[1:0] SYNTHESIZED_WIRE_9;
wire	[1:0] SYNTHESIZED_WIRE_10;
wire	[1:0] SYNTHESIZED_WIRE_11;
wire	[1:0] SYNTHESIZED_WIRE_12;
wire	[1:0] SYNTHESIZED_WIRE_13;
wire	[1:0] SYNTHESIZED_WIRE_14;
wire	[1:0] SYNTHESIZED_WIRE_15;
wire	[1:0] SYNTHESIZED_WIRE_16;
wire	[1:0] SYNTHESIZED_WIRE_17;
wire	[1:0] SYNTHESIZED_WIRE_18;
wire	[1:0] SYNTHESIZED_WIRE_19;
wire	[1:0] SYNTHESIZED_WIRE_20;
wire	[1:0] SYNTHESIZED_WIRE_21;
wire	[1:0] SYNTHESIZED_WIRE_22;
wire	[1:0] SYNTHESIZED_WIRE_23;
wire	[1:0] SYNTHESIZED_WIRE_24;
wire	[1:0] SYNTHESIZED_WIRE_25;
wire	[1:0] SYNTHESIZED_WIRE_26;
wire	[1:0] SYNTHESIZED_WIRE_27;
wire	[1:0] SYNTHESIZED_WIRE_28;
wire	[1:0] SYNTHESIZED_WIRE_29;
wire	[1:0] SYNTHESIZED_WIRE_30;
wire	[1:0] SYNTHESIZED_WIRE_31;
wire	[1:0] SYNTHESIZED_WIRE_32;
wire	[1:0] SYNTHESIZED_WIRE_33;
wire	[1:0] SYNTHESIZED_WIRE_34;
wire	[1:0] SYNTHESIZED_WIRE_35;
wire	[1:0] SYNTHESIZED_WIRE_36;
wire	[1:0] SYNTHESIZED_WIRE_37;
wire	[1:0] SYNTHESIZED_WIRE_38;
wire	[1:0] SYNTHESIZED_WIRE_39;
wire	[1:0] SYNTHESIZED_WIRE_40;
wire	[1:0] SYNTHESIZED_WIRE_41;
wire	[1:0] SYNTHESIZED_WIRE_42;
wire	[1:0] SYNTHESIZED_WIRE_43;
wire	[1:0] SYNTHESIZED_WIRE_44;
wire	[1:0] SYNTHESIZED_WIRE_45;
wire	[1:0] SYNTHESIZED_WIRE_46;
wire	[1:0] SYNTHESIZED_WIRE_47;
wire	[1:0] SYNTHESIZED_WIRE_48;
wire	[1:0] SYNTHESIZED_WIRE_49;
wire	[1:0] SYNTHESIZED_WIRE_50;
wire	[1:0] SYNTHESIZED_WIRE_51;
wire	[1:0] SYNTHESIZED_WIRE_52;
wire	[1:0] SYNTHESIZED_WIRE_53;
wire	[1:0] SYNTHESIZED_WIRE_54;
wire	[1:0] SYNTHESIZED_WIRE_55;
wire	[1:0] SYNTHESIZED_WIRE_56;
wire	[1:0] SYNTHESIZED_WIRE_57;
wire	[1:0] SYNTHESIZED_WIRE_58;
wire	[1:0] SYNTHESIZED_WIRE_59;
wire	[1:0] SYNTHESIZED_WIRE_60;
wire	[1:0] SYNTHESIZED_WIRE_61;
wire	[1:0] SYNTHESIZED_WIRE_62;
wire	[1:0] SYNTHESIZED_WIRE_63;





cvt_128x1_2x64	b2v_inst(
	.Din(tapeData),
	.Dout0_(SYNTHESIZED_WIRE_0),
	.Dout10_(SYNTHESIZED_WIRE_1),
	.Dout11_(SYNTHESIZED_WIRE_2),
	.Dout12_(SYNTHESIZED_WIRE_3),
	.Dout13_(SYNTHESIZED_WIRE_4),
	.Dout14_(SYNTHESIZED_WIRE_5),
	.Dout15_(SYNTHESIZED_WIRE_6),
	.Dout16_(SYNTHESIZED_WIRE_7),
	.Dout17_(SYNTHESIZED_WIRE_8),
	.Dout18_(SYNTHESIZED_WIRE_9),
	.Dout19_(SYNTHESIZED_WIRE_10),
	.Dout1_(SYNTHESIZED_WIRE_11),
	.Dout20_(SYNTHESIZED_WIRE_12),
	.Dout21_(SYNTHESIZED_WIRE_13),
	.Dout22_(SYNTHESIZED_WIRE_14),
	.Dout23_(SYNTHESIZED_WIRE_15),
	.Dout24_(SYNTHESIZED_WIRE_16),
	.Dout25_(SYNTHESIZED_WIRE_17),
	.Dout26_(SYNTHESIZED_WIRE_18),
	.Dout27_(SYNTHESIZED_WIRE_19),
	.Dout28_(SYNTHESIZED_WIRE_20),
	.Dout29_(SYNTHESIZED_WIRE_21),
	.Dout2_(SYNTHESIZED_WIRE_22),
	.Dout30_(SYNTHESIZED_WIRE_23),
	.Dout31_(SYNTHESIZED_WIRE_24),
	.Dout32_(SYNTHESIZED_WIRE_25),
	.Dout33_(SYNTHESIZED_WIRE_26),
	.Dout34_(SYNTHESIZED_WIRE_27),
	.Dout35_(SYNTHESIZED_WIRE_28),
	.Dout36_(SYNTHESIZED_WIRE_29),
	.Dout37_(SYNTHESIZED_WIRE_30),
	.Dout38_(SYNTHESIZED_WIRE_31),
	.Dout39_(SYNTHESIZED_WIRE_32),
	.Dout3_(SYNTHESIZED_WIRE_33),
	.Dout40_(SYNTHESIZED_WIRE_34),
	.Dout41_(SYNTHESIZED_WIRE_35),
	.Dout42_(SYNTHESIZED_WIRE_36),
	.Dout43_(SYNTHESIZED_WIRE_37),
	.Dout44_(SYNTHESIZED_WIRE_38),
	.Dout45_(SYNTHESIZED_WIRE_39),
	.Dout46_(SYNTHESIZED_WIRE_40),
	.Dout47_(SYNTHESIZED_WIRE_41),
	.Dout48_(SYNTHESIZED_WIRE_42),
	.Dout49_(SYNTHESIZED_WIRE_43),
	.Dout4_(SYNTHESIZED_WIRE_44),
	.Dout50_(SYNTHESIZED_WIRE_45),
	.Dout51_(SYNTHESIZED_WIRE_46),
	.Dout52_(SYNTHESIZED_WIRE_47),
	.Dout53_(SYNTHESIZED_WIRE_48),
	.Dout54_(SYNTHESIZED_WIRE_49),
	.Dout55_(SYNTHESIZED_WIRE_50),
	.Dout56_(SYNTHESIZED_WIRE_51),
	.Dout57_(SYNTHESIZED_WIRE_52),
	.Dout58_(SYNTHESIZED_WIRE_53),
	.Dout59_(SYNTHESIZED_WIRE_54),
	.Dout5_(SYNTHESIZED_WIRE_55),
	.Dout60_(SYNTHESIZED_WIRE_56),
	.Dout61_(SYNTHESIZED_WIRE_57),
	.Dout62_(SYNTHESIZED_WIRE_58),
	.Dout63_(SYNTHESIZED_WIRE_59),
	.Dout6_(SYNTHESIZED_WIRE_60),
	.Dout7_(SYNTHESIZED_WIRE_61),
	.Dout8_(SYNTHESIZED_WIRE_62),
	.Dout9_(SYNTHESIZED_WIRE_63));


mux_64x1_2bit	b2v_inst2(
	.Din0_(SYNTHESIZED_WIRE_0),
	.Din10_(SYNTHESIZED_WIRE_1),
	.Din11_(SYNTHESIZED_WIRE_2),
	.Din12_(SYNTHESIZED_WIRE_3),
	.Din13_(SYNTHESIZED_WIRE_4),
	.Din14_(SYNTHESIZED_WIRE_5),
	.Din15_(SYNTHESIZED_WIRE_6),
	.Din16_(SYNTHESIZED_WIRE_7),
	.Din17_(SYNTHESIZED_WIRE_8),
	.Din18_(SYNTHESIZED_WIRE_9),
	.Din19_(SYNTHESIZED_WIRE_10),
	.Din1_(SYNTHESIZED_WIRE_11),
	.Din20_(SYNTHESIZED_WIRE_12),
	.Din21_(SYNTHESIZED_WIRE_13),
	.Din22_(SYNTHESIZED_WIRE_14),
	.Din23_(SYNTHESIZED_WIRE_15),
	.Din24_(SYNTHESIZED_WIRE_16),
	.Din25_(SYNTHESIZED_WIRE_17),
	.Din26_(SYNTHESIZED_WIRE_18),
	.Din27_(SYNTHESIZED_WIRE_19),
	.Din28_(SYNTHESIZED_WIRE_20),
	.Din29_(SYNTHESIZED_WIRE_21),
	.Din2_(SYNTHESIZED_WIRE_22),
	.Din30_(SYNTHESIZED_WIRE_23),
	.Din31_(SYNTHESIZED_WIRE_24),
	.Din32_(SYNTHESIZED_WIRE_25),
	.Din33_(SYNTHESIZED_WIRE_26),
	.Din34_(SYNTHESIZED_WIRE_27),
	.Din35_(SYNTHESIZED_WIRE_28),
	.Din36_(SYNTHESIZED_WIRE_29),
	.Din37_(SYNTHESIZED_WIRE_30),
	.Din38_(SYNTHESIZED_WIRE_31),
	.Din39_(SYNTHESIZED_WIRE_32),
	.Din3_(SYNTHESIZED_WIRE_33),
	.Din40_(SYNTHESIZED_WIRE_34),
	.Din41_(SYNTHESIZED_WIRE_35),
	.Din42_(SYNTHESIZED_WIRE_36),
	.Din43_(SYNTHESIZED_WIRE_37),
	.Din44_(SYNTHESIZED_WIRE_38),
	.Din45_(SYNTHESIZED_WIRE_39),
	.Din46_(SYNTHESIZED_WIRE_40),
	.Din47_(SYNTHESIZED_WIRE_41),
	.Din48_(SYNTHESIZED_WIRE_42),
	.Din49_(SYNTHESIZED_WIRE_43),
	.Din4_(SYNTHESIZED_WIRE_44),
	.Din50_(SYNTHESIZED_WIRE_45),
	.Din51_(SYNTHESIZED_WIRE_46),
	.Din52_(SYNTHESIZED_WIRE_47),
	.Din53_(SYNTHESIZED_WIRE_48),
	.Din54_(SYNTHESIZED_WIRE_49),
	.Din55_(SYNTHESIZED_WIRE_50),
	.Din56_(SYNTHESIZED_WIRE_51),
	.Din57_(SYNTHESIZED_WIRE_52),
	.Din58_(SYNTHESIZED_WIRE_53),
	.Din59_(SYNTHESIZED_WIRE_54),
	.Din5_(SYNTHESIZED_WIRE_55),
	.Din60_(SYNTHESIZED_WIRE_56),
	.Din61_(SYNTHESIZED_WIRE_57),
	.Din62_(SYNTHESIZED_WIRE_58),
	.Din63_(SYNTHESIZED_WIRE_59),
	.Din6_(SYNTHESIZED_WIRE_60),
	.Din7_(SYNTHESIZED_WIRE_61),
	.Din8_(SYNTHESIZED_WIRE_62),
	.Din9_(SYNTHESIZED_WIRE_63),
	.sel(sel),
	.Dout(tapeSymbol));


endmodule
