// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
// CREATED		"Wed Dec 22 01:49:55 2021"

module s8(
	clk,
	rst_n,
	s1,
	resume,
	s8
);


input wire	clk;
input wire	rst_n;
input wire	s1;
input wire	resume;
output reg	s8;

wire	SYNTHESIZED_WIRE_0;





always@(posedge clk or negedge rst_n)
begin
if (!rst_n)
	begin
	s8 <= 0;
	end
else
	begin
	s8 <= SYNTHESIZED_WIRE_0;
	end
end

assign	SYNTHESIZED_WIRE_0 = s1 & resume;


endmodule
