// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
// CREATED		"Tue Dec 21 12:01:21 2021"

module OneHotDecoder2(
	Din,
	Dout
);


input wire	[3:0] Din;
output wire	[1:0] Dout;

wire	[1:0] Dout_ALTERA_SYNTHESIZED;
wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_2;
wire	SYNTHESIZED_WIRE_3;




assign	SYNTHESIZED_WIRE_3 = Din[2] & SYNTHESIZED_WIRE_0;

assign	SYNTHESIZED_WIRE_2 = Din[3] & SYNTHESIZED_WIRE_1;

assign	SYNTHESIZED_WIRE_0 =  ~Din[1];

assign	SYNTHESIZED_WIRE_1 =  ~Din[1];

assign	Dout_ALTERA_SYNTHESIZED[1] = SYNTHESIZED_WIRE_2 | SYNTHESIZED_WIRE_3;

assign	Dout_ALTERA_SYNTHESIZED[0] = Din[3] ^ Din[1];

assign	Dout = Dout_ALTERA_SYNTHESIZED;

endmodule
