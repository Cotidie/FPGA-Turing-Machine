// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition"
// CREATED		"Wed Dec 22 02:12:02 2021"

module triggerMode(
	s,
	mode
);


input wire	[13:0] s;
output wire	[1:0] mode;

wire	[1:0] mode_ALTERA_SYNTHESIZED;




assign	mode_ALTERA_SYNTHESIZED[1] = s[4] | s[2];

assign	mode_ALTERA_SYNTHESIZED[0] = s[4] | s[5] | s[3];

assign	mode = mode_ALTERA_SYNTHESIZED;

endmodule
